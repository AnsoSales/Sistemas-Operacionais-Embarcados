
use IEEE;

entity anso is
	Port();
end;